`define N 256
`define LOG2N 8
